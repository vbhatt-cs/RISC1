library ieee;
use ieee.std_logic_1164.all;
package mem_package is
type ram_t is array (0 to 16383) of std_logic_vector(15 downto 0);
constant MEM_INIT : ram_t := (
0 => "0011001010101011",
1 => "0011010101010100",
2 => "0000010001011000",
3 => "0010010011001001",
4 => "0001011100000010",
5 => "0000100001101000",
6 => "0010011100110010",
7 => "0000110011001000",
8 => "0001001100000001",
9 => "0010100011010001",
10 => "0010001010011000",
11 => "1100001010000011",
12 => "0011101111011101",
13 => "1000010000000100",
14 => "0011001111011101",
15 => "0001000000001011",
16 => "1001010000000000",
17 => "0101101011011110",
18 => "0100110011011110",
19 => "1100101110000010",
20 => "0000010001011000",
21 => "0001100100100000",
22 => "0110100001111111",
23 => "0110000000000000",
24 => "1001011100000000",
25 => "0111110011111111",
others => (others => '0'));
end package mem_package;
